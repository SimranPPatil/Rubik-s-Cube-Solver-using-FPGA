module SRAM_intermediate (input logic Clk, 
				 input logic [15:0] Data_in,
				 output logic [19:0] Data_out,
				 inout wire [15:0] Data  );



endmodule