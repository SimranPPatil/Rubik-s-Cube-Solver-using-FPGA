module ADDER ( input logic Clk, )